**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****

*JSIM model
**HSTP**
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=17ohm, Icrit=0.1mA)
**OPEN**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)
**Low Jc**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.05pF, R0=200ohm, Rn=170ohm, Icrit=10uA)

*** NETLIST FILE ***
**** **** **** **** **** **** **** ****+
*** LIB : ADP_MATSUOKA_LIB
*** CELL: NDROCEX_NEW_VER6TEST
*** VIEW: SCHEMATIC
*** MAY 22 05:01:58 2023
**** **** **** **** **** **** **** ****

*** IJTL
.SUBCKT IJTL          1          2
***       DIN      DOUT
LP2                3         0   0.198PH 
L2                 4         2   1.976PH 
L1                 1         4   4.534PH 
B1                 4         3  JJMOD AREA=2.170
RS1                4         3   5.20OHM *SHUNT=11.30
.ENDS

*** JTL
.SUBCKT JTL          1          2         5
***       DIN      DOUT
R1                 5         6   8.32OHM
LP1                7         0   0.096PH 
LP2                3         0   0.099PH 
L1                 8         9   2.288PH 
L3                 4         2   1.966PH 
L2                 9         4   4.506PH 
LPR1               6         8   0.177PH 
LPIN               1         8   0.317PH 
B1                 9         7  JJMOD AREA=2.160
RS1                9         7   5.23OHM *SHUNT=11.30
B2                 4         3  JJMOD area=2.160
RS2                4         3   5.23OHM *SHUNT=11.30
.ENDS

*** SINK
.SUBCKT SINK          1         5
***       DIN
R2                 4         0   4.08OHM
R1                 5         6   8.32OHM
LP1                7         0   0.130PH 
L1                 8         9   2.272PH 
L2                 9         4   4.766PH 
LPR1               6         8   0.177PH 
LPIN               1         8   0.317PH 
B1                 9         7  jjmod area=2.170
RS1                9         7   5.21OHM *SHUNT=11.30
.ENDS

*** TOP CELL: NDROCEX_NEW_VER6TEST
l1    44    42               2.344pH
l2    42    38               0.670pH
l3    37    38               1.800pH
l4    39    38               1.800pH
l5    32    36               3.851pH
l6    31    35               3.851pH
l7    30    34               1.423pH
l8    31    32               3.851pH
l9    29    33               1.423pH
l10    27    21               3.730pH
l11    26    22               3.730pH
l12    30    27               0.571pH
l13    29    26               0.571pH
l14    21    13               1.990pH
l15    22    15               1.990pH

LP9                0        19   0.184956PH 
LP10               0        24   0.51675PH 
LP11               0        25   0.268894PH 
LP8                0        28   1.25056PH 
LP5               40         0   1.70543PH 
LP4               41         0   2.60469PH 
LP1               43         0   0.289835PH 
LPR1              45        44   0.179528PH 
LPCLK             17        44   0.167969PH 

lX                23         0  10.5PH 
*FIX
lY                20         0  10.312PH 
*FIX
lRST               3         0  12.5PH 
*FIX
lLFB               7         0  31.8062PH 
*FIX


r1    10    45               8.340ohm
*FIX

b1     42    43  jjmod area=1.8     
RS1    42    43               5.381ohm *SHUNT=11.300
*MIN=1.8

b2     37    30  jjmod area=1.77 
RS2    37    30               5.512ohm *SHUNT=11.300

b3     39    29  jjmod area=1.77   
RS3    39    29               5.795ohm *SHUNT=11.300

b4     36    41  jjmod area=2     
RS4    36    41               6.278ohm *SHUNT=11.300

b5     35    40  jjmod area=2     
RS5    35    40               6.278ohm *SHUNT=11.300

b6     32    34  jjmod area=1.000     
RS6    32    34              11.300ohm *SHUNT=11.300
*MIN=1

b7     31    33  jjmod area=1.000     
RS7    31    33              11.300ohm *SHUNT=11.300
*MIN=1

b8     27    28  jjmod area=1.000     
RS8    27    28              11.300ohm *SHUNT=11.300
*MIN=1

b9     26    19  jjmod area=1.000     
RS9    26    19              11.300ohm *SHUNT=11.300
*MIN=1

b10     21    24  jjmod area=1.800     
RS10    21    24               6.647ohm *SHUNT=11.300
*MIN=1.8
*SYN=1

b11     22    25  jjmod area=1.800     
RS11    22    25               6.647ohm *SHUNT=11.300
*MIN=1.8
*SYN=1

K0  LLFB    L7               0.123
K1  LLFB    L8              -0.235
K2  LLFB    L9               0.123

KX    LX    L5              -0.0814
KY    LY    L5              -0.083
KRST  LRST    L6              -0.15


XI13             SINK         14         10
XI10             SINK         16         10
XI33             IJTL         11         12
XI2               JTL         13         14         10
XI3               JTL         15         16         10
XI1               JTL         12         17         10

iBLFB     0     7   PWL(0ps 0mV    50ps                  0.510mA)
*FIX
IINY               0        20  PWL(0PS 0MA 250PS 0MA 251PS 4.12MA 280PS 4.12MA 281PS 0MA 350PS 0MA 351PS 4.12MA 380PS 4.12MA 381PS 0MA)
IINDATA            0        23  PWL(0PS 0MA 350PS 0MA 351PS 1.45MA 380PS 1.45MA 381PS 0MA)
IINRST             0         3  PWL(0PS 0MA 650PS 0MA 651PS 2MA 680PS 2MA 681PS 0MA)

VINCLK            11         0  PULSE(0MV 1.034MV 100PS 1PS 1PS 1PS 100PS)
vB    10     0   PWL(0ps 0mV    50ps                  2.5mV)
*FIX


*** NETLIST FILE ***
.TRAN 0.1ps 1000ps 0ps 1ps

.FILE MARGIN.CSV

.print phase B2
.print phase B3
.print phase B4
.print phase B5
.print phase B8
.print phase B9

.end