**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****

*JSIM model
**HSTP**
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=17ohm, Icrit=0.1mA)
**OPEN**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)
**Low Jc**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.5pF, R0=600ohm, Rn=17ohm, Icrit=0.1mA)


*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : adp_matsuoka_lib
*** Cell: AND_scope
*** View: schematic
*** May 13 18:59:40 2024
**** **** **** **** **** **** **** ****

*** jand
.subckt jand          1          2          3          4        11
***         a         b         c       clk
r3                11        12  33.52ohm
r8                11        13   8.32ohm 
*FIX
r1                11        14  17.52ohm
r5                11        15   8.32ohm 
*FIX
r4                11        16  14.88ohm
r2                11        17  17.52ohm
r6                11        18   8.32ohm 
*FIX

l1                26        27   2.844pH fcheck 
l2                52        53   2.904pH fcheck 
l3                44        33   2.054pH fcheck 
l4                47        42   2.057pH fcheck 
l5                31        32   2.132pH fcheck 
l6                31        41   2.171pH fcheck 
l7                36        37   1.924pH fcheck 
l8                23        21   0.039pH fcheck 
l9                21        20   2.600pH fcheck 
l10               20         3   2.470pH fcheck 
l11               43        44   5.075pH fcheck 
l12               46        47   4.800pH fcheck 
l13               28        43   2.389pH fcheck 
l14               50        46   2.410pH fcheck 
l15               33        25   9.521pH fcheck 
l16               42        51   9.547pH fcheck 
l17               29        30   2.192pH fcheck 
l18               30        39   5.021pH fcheck 
l19               39        36   0.239pH fcheck 
l20               22        23   0.499pH fcheck 
l21               25        26   0.148pH fcheck 
l22               51        52   0.179pH fcheck 
l23               37        31   0.010pH fcheck 




LP1               19         0   0.255pH fcheck 
LPR3              12        21   1.901pH fcheck 
LP9               24         0   0.174pH fcheck 
LPR5              15        28   0.166pH fcheck 
LPCLK              4        29   0.291pH fcheck 
LPR8              13        29   0.166pH fcheck 
LPR1              14        33   0.013pH fcheck 
LP7               34         0   0.299pH fcheck 
LP12              35         0   0.203pH fcheck 
LP15              38         0   0.190pH fcheck 
LP14              40         0   0.187pH fcheck 
LPR4              16        36   0.850pH fcheck 
LPR2              17        42   0.010pH fcheck 
LP13              45         0   0.195pH fcheck 
LP11              48         0   0.203pH fcheck 
LP10              49         0   0.221pH fcheck 
LPA                1        28   0.291pH fcheck 
LPB                2        50   0.286pH fcheck 
LPR6              18        50   0.172pH fcheck 
LP8               54         0   0.211pH fcheck 
LP2               55         0   0.229pH fcheck 

b1                25        19  jjmod area=1.21
RS1               25        19   9.34ohm *SHUNT=11.30
b2                51        55  jjmod area=1.21
RS2               51        55   9.34ohm *SHUNT=11.30
b3                26        32  jjmod area=1.05
RS3               26        32  10.76ohm *SHUNT=11.30
b4                52        41  jjmod area=1.05
RS4               52        41  10.76ohm *SHUNT=11.30
b5                27        22  jjmod area=1.38
RS5               27        22   8.19ohm *SHUNT=11.30
b6                53        22  jjmod area=1.38
RS6               53        22   8.19ohm *SHUNT=11.30
b7                23        34  jjmod area=1.56
RS7               23        34   7.23ohm *SHUNT=11.30
Bb                37        54  jjmod area=1.38
RS8               37        54   8.19ohm *SHUNT=11.30
b9                20        24  jjmod area=2.61
RS9               20        24   4.33ohm *SHUNT=11.30
*FIX
b10               44        49  jjmod area=1.75
RS10              44        49   6.44ohm *SHUNT=11.30
b11               47        48  jjmod area=1.75
RS11              47        48   6.44ohm *SHUNT=11.30
b12               43        35  jjmod area=2.17
RS12              43        35   5.20ohm *SHUNT=11.30
*FIX
b13               46        45  jjmod area=2.17
RS13              46        45   5.20ohm *SHUNT=11.30
*FIX
b14               39        40  jjmod area=1.26
RS14              39        40   8.93ohm *SHUNT=11.30
b15               30        38  jjmod area=2.17
RS15              30        38   5.20ohm *SHUNT=11.30
*FIX
.ends

*** jtl
.subckt jtl         56         57        17
***       din      dout
B1                53        58  jjmod area=2.16
RS1               53        58   5.23ohm *SHUNT=11.30
B2                22        27  jjmod area=2.16
RS2               22        27   5.23ohm *SHUNT=11.30
LP1               58         0   0.096pH fcheck 
LP2               27         0   0.099pH fcheck 
L1                44        53   2.288pH fcheck 
L3                22        57   1.963pH fcheck 
L2                53        22   4.506pH fcheck 
LPR1              13        44   0.177pH fcheck 
LPIN              56        44   0.317pH fcheck 
R1                17        13   8.32ohm
.ends

*** ijtl
.subckt ijtl         56         57
***       din      dout
B1                39        50  jjmod area=2.17
RS1               39        50   5.20ohm *SHUNT=11.30
LP2               50         0   0.198pH fcheck 
L2                39        57   1.976pH fcheck 
L1                56        39   4.534pH fcheck 
.ends

*** sink
.subckt sink         56        58
***       din
B1                31        28  jjmod area=2.17
RS1               31        28   5.21ohm *SHUNT=11.30
LP1               28         0   0.130pH fcheck 
L1                46        31   2.272pH fcheck 
L2                31        42   4.766pH fcheck 
LPR1              53        46   0.177pH fcheck 
LPIN              56        46   0.317pH fcheck 
R2                42         0   4.08ohm
R1                58        53   8.32ohm
.ends

*** top cell: AND_scope
XI0              jand         39         43         44         42         29
XI7               jtl         44         47         29
XI4               jtl         36         43         29
XI2               jtl         46         39         29
XI6               jtl         37         42         29
XI5              ijtl         59         37
XI3              ijtl         60         36
XI1              ijtl         61         46
XI8              sink         47         29


vb                29         0  PWL(0ps 0mv 50ps 2.5mv) 
*FIX
Vinclk            59         0  PULSE(0mv 1.034mv 100ps 1ps 1ps 1ps 100ps)

Vina              61         0  PWL(0ps 0mv 150ps 0mv 151ps 2.068mv 152ps 0mv 320ps 0mv 321ps 2.068mv 322ps 0mv 520ps 0mv 521ps 2.068mv 522ps 0mv 570ps 0mv 571ps 2.068mv 572ps 0mv)
Vinb              60         0  PWL(0ps 0mv 250ps 0mv 251ps 2.068mv 252ps 0mv 370ps 0mv 371ps 2.068mv 372ps 0mv 620ps 0mv 621ps 2.068mv 622ps 0mv 670ps 0mv 671ps 2.068mv 672ps 0mv)




*** netlist file ***

*** jsim input file ***

*** jsim input file ***
.tran 1ps 800ps 0ps 0.2ps:
.file a.csv

.print phase XI0_B1
.print phase XI0_B2
.print phase XI0_B3
.print phase XI0_B4
.print phase XI0_B7



.end