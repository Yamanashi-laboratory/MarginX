**** **** **** **** **** **** **** **** **** **** **** 
*JSIM CONTROL FILE FOR CADENCE BY KAMEDA@CQ.JP.NEC.COM
**** **** **** **** **** **** **** **** **** **** ****

*JSIM MODEL
.MODEL JJMOD JJ(RTYPE=1, VG=2.8MV, CAP=0.064PF, R0=100OHM, RN=16OHM, ICRIT=0.1MA)

*** NETLIST FILE ***
**** **** **** **** **** **** **** ****+
*** LIB : ADP_KUNIHIRO_LIB
*** CELL: TEST_DFF
*** VIEW: SCHEMATIC
*** FEB 10 21:27:58 2022
**** **** **** **** **** **** **** ****

*** IJTL
.SUBCKT IJTL          1          2
***       DIN      DOUT
LP2                3         0   0.198PH FCHECK
L2                 4         2   1.976PH FCHECK
L1                 1         4   4.534PH FCHECK
B1                 4         3  JJMOD AREA=2.170
RS1                4         3   5.20OHM *SHUNT=11.30
.ENDS

*** JTL
.SUBCKT JTL          1          2         5
***       DIN      DOUT
R1                 5         6   8.32OHM
LP1                7         0   0.096PH FCHECK
LP2                3         0   0.099PH FCHECK
L1                 8         9   2.288PH FCHECK
L3                 4         2   1.963PH FCHECK
L2                 9         4   4.506PH FCHECK
LPR1               6         8   0.177PH FCHECK
LPIN               1         8   0.317PH FCHECK
B1                 9         7  JJMOD AREA=2.160
RS1                9         7   5.23OHM *SHUNT=11.30
B2                 4         3  JJMOD AREA=2.160
RS2                4         3   5.23OHM *SHUNT=11.30
.ENDS

*** OPT_DFF
.SUBCKT OPT_DFF         10          1          2        29
***       CLK       DIN      DOUT
b6                18         7  JJMOD AREA=2.160
RS6 18 7 5.231OHM
*FIX
b5                11         4  JJMOD AREA=2.160
RS5 11 4 5.231OHM
*FIX
b4                19        20  JJMOD AREA=1.839
RS4 19 20 6.146OHM
b3                14        15  JJMOD AREA=1.746
RS3 14 15 6.472OHM
b2                12        13  JJMOD AREA=2.160
RS2 12 13 5.231OHM
*FIX

b1                16        17  JJMOD AREA=1.799
RS1 16 17 6.281OHM

LPR3              22        21   0.159PH FCHECK
LPR2              26        25   0.156PH FCHECK
LPR1              23        24   0.104PH FCHECK
LPCLK             10        21   0.361PH FCHECK
LP6                7         0   0.127PH FCHECK
LP5                4         0   0.096PH FCHECK
LP4               20         0   0.276PH FCHECK
LP3               15         0   0.104PH FCHECK
LP2               13         0   0.094PH FCHECK
LPIN               1        25   0.328PH FCHECK
L9                16        19   0.042PH FCHECK
l8 18 2 2.591PH FCHECK
l7 25 12 2.903PH FCHECK
l6 21 11 2.354PH FCHECK
l5 12 14 3.608PH FCHECK
l4 19 18 3.786PH FCHECK
l3 24 16 4.132PH FCHECK
l2 14 24 2.083PH FCHECK
l1 11 17 3.654PH FCHECK
r3 29 22 8.320OHM
r2 29 26 8.320OHM
r1 29 23 11.441OHM
.ENDS

*** SINK
.SUBCKT SINK          1         5
***       DIN
R2                 4         0   4.08OHM
R1                 5         6   8.32OHM
LP1                7         0   0.130PH FCHECK
L1                 8         9   2.272PH FCHECK
L2                 9         4   4.766PH FCHECK
LPR1               6         8   0.177PH FCHECK
LPIN               1         8   0.317PH FCHECK
B1                 9         7  JJMOD AREA=2.170
RS1                9         7   5.21OHM *SHUNT=11.30
.ENDS

*** TOP CELL: TEST_DFF
VINCLK            30         0  PWL(0PS 0MV 100PS 0MV 101PS 1.035MV 102PS 1.035MV 103PS 0MV 300PS 0MV 301PS 1.035MV 302PS 1.035MV 303PS 0MV 400PS 0MV 401PS 1.035MV 402PS 1.035MV 403PS 0MV 600PS 0MV 601PS 1.035MV 602PS 1.035MV 603PS 0MV)
VINDIN               31         0  PWL(0PS 0MV 200PS 0MV 201PS 1.035MV 202PS 1.035MV 203PS 0MV 500PS 0MV 501PS 1.035MV 502PS 1.035MV 503PS 0MV)
vb 32 0 PWL(0PS 0MV 20PS 2.5MV)
*FIX
XI1              IJTL         30         33
XI3              IJTL         31         34
XI2               JTL         33          9         32
XI6               JTL         35         36         32
XI4               JTL         34         37         32
XI5           OPT_DFF          9         37         35         32
XI7              SINK         36         32


*** netlist file ***
.TRAN 0.1ps 750ps 0ps 1ps
.FILE si_dff.csv
.print phase B1.XI1
.print phase B1.XI3
.print phase B1.XI7



.end
