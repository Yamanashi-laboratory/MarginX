**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****

*JSIM model
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)

*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : nec_nakaishi_lib
*** Cell: NDRO
*** View: schematic
*** Nov 16 15:28:27 2017
**** **** **** **** **** **** **** ****

*** top cell: NDRO
B25                1         2  jjmod area=2.16
RS25               1         2   1.73ohm *SHUNT=3.73
B22                3         4  jjmod area=2.16
RS22               3         4   1.73ohm *SHUNT=3.73
B21                5         6  jjmod area=2.16
RS21               5         6   1.73ohm *SHUNT=3.73
B20                7         8  jjmod area=2.16
RS20               7         8   1.73ohm *SHUNT=3.73
B19                9        10  jjmod area=2.16
RS19               9        10   1.73ohm *SHUNT=3.73
B18               11        12  jjmod area=2.16
RS18              11        12   1.73ohm *SHUNT=3.73
B17               13        14  jjmod area=2.16
RS17              13        14   1.73ohm *SHUNT=3.73
B23               15        16  jjmod area=2.16
RS23              15        16   1.73ohm *SHUNT=3.73
B16               17        18  jjmod area=2.16
RS16              17        18   1.73ohm *SHUNT=3.73
B15               19        20  jjmod area=2.16
RS15              19        20   1.73ohm *SHUNT=3.73
B14               21        22  jjmod area=2.16  
RS14              21        22   1.73ohm *SHUNT=3.73
B13               23        24  jjmod area=2.16
RS13              23        24   1.73ohm *SHUNT=3.73
B12               25        26  jjmod area=2.16
RS12              25        26   1.73ohm *SHUNT=3.73
B0                27        28  jjmod area=2.16
RS0               27        28   1.73ohm *SHUNT=3.73
b10     29    30  jjmod area=1.933     
RS10    29    30               1.929ohm *SHUNT=3.730
b11     31    32  jjmod area=2.237     
RS11    31    32               1.667ohm *SHUNT=3.730
b5     33    34  jjmod area=2.621     
RS5    33    34               1.423ohm *SHUNT=3.730
b7     35    36  jjmod area=2.246     
RS7    35    36               1.661ohm *SHUNT=3.730
b8     36    37  jjmod area=1.456     
RS8    36    37               2.562ohm *SHUNT=3.730
b4     38    33  jjmod area=2.464     
RS4    38    33               1.514ohm *SHUNT=3.730
b9     39    40  jjmod area=1.107     
RS9    39    40               3.370ohm *SHUNT=3.730
B24               41        42  jjmod area=2.16
RS24              41        42   1.73ohm *SHUNT=3.73
b3     43    44  jjmod area=2.409     
RS3    43    44               1.548ohm *SHUNT=3.730
b6     45    46  jjmod area=2.398     
RS6    45    46               1.556ohm *SHUNT=3.730
b1     47    48  jjmod area=2.318     
RS1    47    48               1.609ohm *SHUNT=3.730

b2     47    49  jjmod area=2.180     
RS2    47    49               1.711ohm *SHUNT=3.730
***mid = 1.641

L64                2         0   0.205pH fcheck
L63                1        50   1.890pH fcheck
L62               51         1   4.945pH fcheck
L61               52        41   4.945pH fcheck
L56               53        15   4.945pH fcheck
L55               54        55   0.359pH fcheck
L54               56        55   0.270pH fcheck
L53               55         5   2.379pH fcheck
L52                4         0   0.234pH fcheck
L51                6         0   0.250pH fcheck
L50                5         3   5.130pH fcheck
L49               57         7   4.945pH fcheck
L48               58        57   4.277pH fcheck
L47                3        57   0.091pH fcheck
L46                7        59   5.000pH fcheck
L45                8         0   0.205pH fcheck
L59               42         0   0.205pH fcheck
L44               10         0   0.205pH fcheck
L43                9        60   1.890pH fcheck
L42               13        61   0.091pH fcheck
L41               62        61   4.277pH fcheck
L40               61         9   4.945pH fcheck
L39               11        13   5.130pH fcheck
L38               12         0   0.250pH fcheck
L37               14         0   0.234pH fcheck
L36               63        11   2.379pH fcheck
L35               64        63   0.270pH fcheck
L34               65        63   0.359pH fcheck
L33               66        67   0.359pH fcheck
L32               68        67   0.270pH fcheck
L31               67        19   2.379pH fcheck
L30               18         0   0.234pH fcheck
L29               20         0   0.250pH fcheck
L28               19        17   5.130pH fcheck
L27               69        21   4.945pH fcheck
L26               70        69   4.277pH fcheck
L25               17        69   0.091pH fcheck
L24               21        71   1.890pH fcheck
L23               22         0   0.205pH fcheck
L57               15        65   1.890pH fcheck
L22               24         0   0.205pH fcheck
L21               23        72   1.890pH fcheck
L20               27        73   0.091pH fcheck
L19               74        73   4.277pH fcheck
L18               73        23   4.945pH fcheck
L17               25        27   5.130pH fcheck
L16               26         0   0.250pH fcheck
LP2               28         0   0.234pH fcheck
L15               75        25   2.379pH fcheck
L0                76        75   0.270pH fcheck
LPIN              50        75   0.359pH fcheck
L60               41        66   1.890pH fcheck
l11    29    31               4.791pH
LP10              30         0   0.112pH fcheck
LP11              32         0   0.120pH fcheck
L12               31        54   2.096pH fcheck
l2    49    77               2.639pH
LP8               37         0   0.255pH fcheck
l14    36    78               0.784pH
l8    33    39               2.584pH
LP5               34         0   0.268pH fcheck
l13    77    29               0.806pH
l9    40    79               0.399pH
l10    79    77               0.396pH
l7    78    39               3.173pH
LPR5              80        79   0.205pH fcheck
LPR4              81        78   0.328pH fcheck
L58               16         0   0.205pH fcheck
LPR3              82        83   0.244pH fcheck
L5                83        45   2.205pH fcheck
LPDIN             72        83   0.234pH fcheck
LPR2              84        85   0.237pH fcheck
LPRESET           71        85   0.200pH fcheck
L3                85        43   2.527pH fcheck
LPCLK             60        86   0.203pH fcheck
LPR1              87        86   0.239pH fcheck
L1                86        47   2.137pH fcheck
LP6               46         0   0.112pH fcheck
l6    45    35               3.535pH
l4    43    38               2.594pH
LP3               44         0   0.156pH fcheck
LP1               48         0   0.177pH fcheck
R16               59         0   10.00ohm
R12               98        56   8.34ohm
R11               98        58  16.65ohm
R10               98        62  16.65ohm
R9                98        64   8.34ohm
R8                98        68   8.34ohm
R7                98        70  16.65ohm
R6                98        74  16.65ohm
R0                98        76   8.34ohm
r5    80    98              30.039ohm
r4    98    81              31.565ohm
R2                98        84   8.34ohm
R3                98        82   8.34ohm
R1                98        87   8.34ohm


V0                51         0  PWL(0ps 0mV 550ps 0mV 552ps 1.034mV 554ps 0mV 650ps 0mV 652ps 1.034mV 654ps 0mV 950ps 0mV 952ps 1.034mV 954ps 0mV)
V1                52         0  PWL(0ps 0mV 750ps 0mV 752ps 1.034mV 754ps 0mV 850ps 0mV 852ps 1.034mV 854ps 0mV)
V2                53         0  PWL(0ps 0mV 500ps 0mV 502ps 1.034mV 504ps 0mV 600ps 0mV 602ps 1.034mV 604ps 0mV 700ps 0mV 702ps 1.034mV 704ps 0mV 800ps 0mV 802ps 1.034mV 804ps 0mV 900ps 0mV 902ps 1.034mV 904ps 0mV 1000ps 0mV 1002ps 1.034mV 1004ps 0mV 1100ps 0mV 1102ps 1.034mV 1104ps 0mV)

vb    98     0   PWL(0ps 0mV    20ps                  2.500mV)
*FIX
.tran 0.1ps 1.2ns 0.4ns 0.2ps
 

.FILE ex03_out.CSV

.print phase B11
.print phase B7
.print phase B4
.print phase B2
.print phase B9


*** netlist file ***

*** jsim input file ***

*** jsim input file ***
