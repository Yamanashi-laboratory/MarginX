**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****

*JSIM model
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=16ohm, Icrit=0.1mA)

*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : adp_kunihiro_lib
*** Cell: test_dff
*** View: schematic
*** Feb 10 21:27:58 2022
**** **** **** **** **** **** **** ****

*** ijtl
.subckt ijtl          1          2
***       din      dout
LP2                3         0   0.198pH fcheck
L2                 4         2   1.976pH fcheck
L1                 1         4   4.534pH fcheck
B1                 4         3  jjmod area=2.17
RS1                4         3   5.20ohm *SHUNT=11.30
.ends

*** jtl
.subckt jtl          1          2         5
***       din      dout
R1                 5         6   8.32ohm
LP1                7         0   0.096pH fcheck
LP2                3         0   0.099pH fcheck
L1                 8         9   2.288pH fcheck
L3                 4         2   1.963pH fcheck
L2                 9         4   4.506pH fcheck
LPR1               6         8   0.177pH fcheck
LPIN               1         8   0.317pH fcheck
B1                 9         7  jjmod area=2.16
RS1                9         7   5.23ohm *SHUNT=11.30
B2                 4         3  jjmod area=2.16
RS2                4         3   5.23ohm *SHUNT=11.30
.ends

*** opt_dff
.subckt opt_dff         10          1          2        29
***       clk       din      dout
b6     18     7  jjmod area=2.659     
RS6    18     7               4.249ohm *SHUNT=11.300
b5     11     4  jjmod area=1.321     
RS5    11     4               8.556ohm *SHUNT=11.300
b4     19    20  jjmod area=1.374     
RS4    19    20               8.227ohm *SHUNT=11.300
b3     14    15  jjmod area=1.644     
RS3    14    15               6.875ohm *SHUNT=11.300
b2     12    13  jjmod area=1.208     
RS2    12    13               9.356ohm *SHUNT=11.300
b1     16    17  jjmod area=1.598     
RS1    16    17               7.071ohm *SHUNT=11.300
LPR3              22        21   0.159pH fcheck
LPR2              26        25   0.156pH fcheck
LPR1              23        24   0.104pH fcheck
LPCLK             10        21   0.361pH fcheck
LP6                7         0   0.127pH fcheck
LP5                4         0   0.096pH fcheck
LP4               20         0   0.276pH fcheck
LP3               15         0   0.104pH fcheck
LP2               13         0   0.094pH fcheck
LPIN               1        25   0.328pH fcheck
L9                16        19   0.042pH fcheck
l8    18     2               1.531pH
l7    25    12               2.322pH
l6    21    11               1.848pH
l5    12    14               2.954pH
l4    19    18               4.006pH
l3    24    16               5.887pH
l2    14    24               1.265pH
l1    11    17               2.208pH
r3    29    22              18.533ohm
r2    29    26              16.111ohm
r1    29    23              40.969ohm
.ends

*** sink
.subckt sink          1         5
***       din
R2                 4         0   4.08ohm
R1                 5         6   8.32ohm
LP1                7         0   0.130pH fcheck
L1                 8         9   2.272pH fcheck
L2                 9         4   4.766pH fcheck
LPR1               6         8   0.177pH fcheck
LPIN               1         8   0.317pH fcheck
B1                 9         7  jjmod area=2.17
RS1                9         7   5.21ohm *SHUNT=11.30
.ends

*** top cell: test_dff
Vinclk            30         0  PWL(0ps 0mv 100ps 0mv 101ps 1.035mv 102ps 1.035mv 103ps 0mv 300ps 0mv 301ps 1.035mv 302ps 1.035mv 303ps 0mv 400ps 0mv 401ps 1.035mv 402ps 1.035mv 403ps 0mv 600ps 0mv 601ps 1.035mv 602ps 1.035mv 603ps 0mv)
Vindin               31         0  PWL(0ps 0mv 200ps 0mv 201ps 1.035mv 202ps 1.035mv 203ps 0mv 500ps 0mv 501ps 1.035mv 502ps 1.035mv 503ps 0mv)
vb    32     0   PWL(0ps 0mV    20ps                  2.500mV)
*FIX
XI1              ijtl         30         33
XI3              ijtl         31         34
XI2               jtl         33          9         32
XI6               jtl         35         36         32
XI4               jtl         34         37         32
XI5           opt_dff          9         37         35         32
XI7              sink         36         32

*** netlist file ***
.tran 0.1ps 750ps 0ps 1ps
.FILE ./test/dff_out.CSV

.print phase B1.XI5
.print phase B3.XI5
.print phase B4.XI5

*** jsim input file ***

*** jsim input file ***
