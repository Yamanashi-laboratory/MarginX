**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****

*JSIM model
**HSTP**
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=17ohm, Icrit=0.1mA)
**OPEN**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)
**Low Jc**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.05pF, R0=200ohm, Rn=170ohm, Icrit=10uA)


*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : hstp_yahata_lib
*** Cell: test_ORC_ver3x1
*** View: schematic
*** Jul 17 11:16:49 2023
**** **** **** **** **** **** **** ****



*** ijtl
.subckt ijtl         50         51
***       din      dout
L1                50        52   4.776pH fcheck
L3                52        51   1.620pH fcheck
LP1               16         0   0.218pH fcheck
B1                52        16  jjmod area=2.13
RS1               52        16   5.31ohm *SHUNT=11.30
.ends

*** jtl
.subckt jtl         50         51        53
***       din      dout
R1                53        54   8.32ohm
LPIN              50        55   0.840pH fcheck
LPR1              54        55   3.588pH fcheck
L2                11        21   4.776pH fcheck
L3                21        51   1.620pH fcheck
L1                55        11   2.467pH fcheck
LP2               16         0   0.218pH fcheck
LP1               14         0   0.224pH fcheck
B2                21        16  jjmod area=2.13
RS2               21        16   5.31ohm *SHUNT=11.30
B1                11        14  jjmod area=2.13
RS1               11        14   5.31ohm *SHUNT=11.30
.ends

*** sink
.subckt sink         50        17
***       din
R1                17        56   8.32ohm
R2                12         0   4.02ohm
LPIN              50        57   0.840pH fcheck
LPR1              56        57   3.588pH fcheck
L3                14        12   4.792pH fcheck
L1                57        14   2.475pH fcheck
LP1               21         0   0.218pH fcheck
B1                14        21  jjmod area=2.13
RS1               14        21   5.31ohm *SHUNT=11.30
.ends

*** ORC_ver3x1
.subckt ORC_ver3x1          1          2          3          4          5        49
***         a         b         c     c_bar       clk
***����L2���߂��l���Ƃ�����L5
l1                44        42   3.301pH fcheck 
l2                39        32   3.301pH fcheck 
l3                36        34   3.301pH fcheck 
L4                42        30   3.301pH fcheck 
L5                32        17   1.000pH fcheck 
L6                34        29   3.301pH fcheck 
L7                30        31   1.481pH fcheck
L8                28        29   1.481pH fcheck 
L9                27        24   0.513pH fcheck 
L10               17        19   1.955pH fcheck 
L11               24        25   3.300pH fcheck 
L12               17        18   1.588pH fcheck 
L13               22        21   4.547pH fcheck 
l14               16        20   3.223pH fcheck 
L15               21        11   2.306pH fcheck 
L16               16        14   0.825pH fcheck 
L17               11         9   0.471pH fcheck 
L18               14        12   5.000pH fcheck 
L19                9         7   4.042pH fcheck 
L20               12         4   2.003pH fcheck 
L21                7         3   2.004pH fcheck 
l22                6         0  29.162pH fcheck 

LPR1              44        45   4.831pH fcheck 
LPR2              39        40   5.061pH fcheck 
LPR3              36        37   4.831pH fcheck 
LPR4              24        26   3.500pH fcheck 



LPA                1        44   0.842pH fcheck 
LPCLK              5        39   0.842pH fcheck 
LPB                2        36   0.842pH fcheck 


LP1               43         0   0.200pH fcheck
LP2               38         0   0.200pH fcheck
LP3               35         0   0.200pH fcheck
LP4               41         0   0.200pH fcheck
LP5               33         0   0.200pH fcheck
LP11              23         0   0.200pH fcheck
LP14              10         0   0.200pH fcheck
LP13              15         0   0.200pH fcheck
LP15              13         0   0.200pH fcheck
LP16               8         0   0.200pH fcheck


r1                45        49   8.32ohm 
r2                40        49   7.44ohm 
r3                37        49   8.32ohm 
r4                26        49   9.60ohm 

b1                42        43  jjmod area=2.13 
RS1               42        43   5.30ohm *SHUNT=11.30
b2                32        38  jjmod area=2.13 
RS2               32        38   5.30ohm *SHUNT=11.30
b3                34        35  jjmod area=2.13 
RS3               34        35   5.30ohm *SHUNT=11.30
b4                30        41  jjmod area=2.13 
RS4               30        41   5.30ohm *SHUNT=11.30
b5                29        33  jjmod area=2.13 
RS5               29        33   5.30ohm *SHUNT=11.30
b6                31        27  jjmod area=1.80 
RS6               31        27   6.29ohm *SHUNT=11.30
b7                28        27  jjmod area=1.80 
RS7               28        27   6.29ohm *SHUNT=11.30
b8                19        16  jjmod area=1 
RS8               19        16  11.30ohm *SHUNT=11.30
b9                25        22  jjmod area=2.07 
RS9               25        22   5.45ohm *SHUNT=11.30
b10               18        11  jjmod area=1.5 
RS10              18        11   11.30ohm *SHUNT=11.30
b11               22        23  jjmod area=2.02 
RS11              22        23   5.61ohm *SHUNT=11.30
b12               21        20  jjmod area=0.8 
RS12              21        20  13.95ohm *SHUNT=11.30
b13               14        15  jjmod area=0.71 
RS13              14        15  16.01ohm *SHUNT=11.30
b14                9        10  jjmod area=1.05 
RS14               9        10  10.76ohm *SHUNT=11.30
b15               12        13  jjmod area=1.00 
RS15              12        13  11.30ohm *SHUNT=11.30
b16                7         8  jjmod area=1.25 
RS16               7         8   9.01ohm *SHUNT=11.30


k2                L13        L22 0.227 
k1                L14        L22 0.245
ib                 0         6  PWL(0ps 0mA 50ps 0.5mA) 


.ends

*** top cell: test_ORC_ver3x1
XI0        ORC_ver3x1         56         14         39         32         58         42
vb                42         0  PWL(0ps 0mV 50ps 2.5mV) 

Vinclk            24         0  PWL(0ps 0mv 200ps 0mV 201ps 1.034mV 202ps 1.034mV 203ps 0mV 400ps 0mV 401ps 1.034mV 402ps 1.034mV 403ps 0mV 600ps 0mV 601ps 1.034mV 602ps 1.034mV 603ps 0mV 800ps 0mV 801ps 1.034mV 802ps 1.034mV 803ps 0mV)
Vina              11         0  PWL(0ps 0mv 250ps 0mV 251ps 1.034mV 252ps 1.034mV 253ps 0mV 350ps 0mV 351ps 1.034mV 352ps 1.034mV 353ps 0mV 650ps 0mV 651ps 1.034mV 652ps 1.034mV 653ps 0mV 750ps 0mV 751ps 1.034mV 752ps 1.034mV 753ps 0mV)
Vinb              30         0  PWL(0ps 0mv 450ps 0mV 451ps 1.034mV 452ps 1.034mV 453ps 0mV 550ps 0mV 551ps 1.034mV 552ps 1.034mV 553ps 0mV 650ps 0mV 651ps 1.034mV 652ps 1.034mV 653ps 0mV 750ps 0mV 751ps 1.034mV 752ps 1.034mV 753ps 0mV)


Xijtlb           ijtl         30         17
Xijtlclk         ijtl         24         27
Xijtla           ijtl         11         22
Xjtlc2            jtl         36         21         42
Xjtlcbar2         jtl         44         16         42
Xjtlc1            jtl         39         36         42
Xjtlcbar1         jtl         32         44         42
Xjtlb2            jtl          9         14         42
Xjtlclk2          jtl         12         58         42
Xjtla2            jtl         59         56         42
Xjtlb1            jtl         17          9         42
Xjtlclk1          jtl         27         12         42
Xjtla1            jtl         22         59         42
Xsinkc           sink         21         42
Xsinkcbar        sink         16         42


.tran 0.1ps 1000ps 0ps 1ps
.FILE MARGIN.txt

.print phase B6.XI0
.print phase B7.XI0
.print phase B8.XI0
.print phase B9.XI0
.print phase B10.XI0
.print phase B11.XI0
.print phase B12.XI0
.print phase B13.XI0
.print phase B14.XI0
.end

