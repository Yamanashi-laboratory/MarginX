**** **** **** **** **** **** **** **** **** **** **** 
*JSIM control file for CADENCE by kameda@cq.jp.nec.com
**** **** **** **** **** **** **** **** **** **** ****
*BIN=1
*JSIM model
**HSTP**
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=17ohm, Icrit=0.1mA)
**OPEN**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)
**Low Jc**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.5pF, R0=600ohm, Rn=17ohm, Icrit=0.1mA)


*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : adp_matsuoka_lib
*** Cell: ndrotest
*** View: schematic
*** Apr 12 02:42:34 2024
**** **** **** **** **** **** **** ****

*** ijtl
.subckt ijtl          1          2
***       din      dout
B1                 3         4  jjmod area=2.17
RS1                3         4   5.20ohm *SHUNT=11.30
LP2                4         0   0.198pH fcheck
L2                 3         2   1.976pH fcheck
L1                 1         3   4.534pH fcheck
.ends

*** jtl
.subckt jtl          1          2        11
***       din      dout
B1                 5         6  jjmod area=2.16
RS1                5         6   5.23ohm *SHUNT=11.30
B2                 7         8  jjmod area=2.16
RS2                7         8   5.23ohm *SHUNT=11.30
LP1                6         0   0.096pH fcheck
LP2                8         0   0.099pH fcheck
L1                 9         5   2.288pH fcheck
L3                 7         2   1.963pH fcheck
L2                 5         7   4.506pH fcheck
LPR1              10         9   0.177pH fcheck
LPIN               1         9   0.317pH fcheck
R1                11        10   8.32ohm
.ends

*** sink
.subckt sink          1         6
***       din
B1                12        13  jjmod area=2.17
RS1               12        13   5.21ohm *SHUNT=11.30
LP1               13         0   0.130pH fcheck
L1                14        12   2.272pH fcheck
L2                12        15   4.766pH fcheck
LPR1               5        14   0.177pH fcheck
LPIN               1        14   0.317pH fcheck
R2                15         0   4.08ohm
R1                 6         5   8.32ohm
.ends

*** top cell: ndrotest
l1    53    54               2.074pH
l2    45    36               2.840pH
l3    55    46               2.355pH
l4    46    47               2.712pH
l5    56    48               2.255pH
l6    48    49               3.734pH
l7    40    38               3.481pH
l8    41    40               3.206pH
l9    39    34               0.471pH
l10    34    36               0.397pH
l11    32    30               5.145pH
l12    30    22               1.707pH
l13    36    32               0.924pH
l14    42    38               0.803pH

LP11              31         0   0.133pH fcheck
LPR5              33        34   0.070pH fcheck
LP10              35         0   0.151pH fcheck
LPR4              37        38   0.434pH fcheck
LP5               43         0   0.159pH fcheck
LP8               44         0   0.172pH fcheck
LP1               50         0   0.146pH fcheck
LP3               51         0   0.148pH fcheck
LP6               52         0   0.127pH fcheck
LPR1              57        53   0.198pH fcheck
LPR2              58        55   0.198pH fcheck
LPR3              59        56   0.200pH fcheck
LPCLK             24        53   0.216pH fcheck
LPDIN             14        56   0.237pH fcheck
LPRESET           23        55   0.216pH fcheck

r1     4    57               8.340ohm
*FIX
r2     4    58               8.340ohm
*FIX
r3     4    59               8.340ohm
*FIX

r4     4    37              24.313ohm
r5    33     4              22.475ohm

b1    54    50  jjmod area=2.100     
RS1    54    50               5.381ohm  *SHUNT=11.300
*FIX
b2    54    45  jjmod area=1.535     
RS2    54    45               7.360ohm  *SHUNT=11.300
b3    46    51  jjmod area=2.180     
RS3    46    51               5.183ohm  *SHUNT=11.300
*FIX
b4    47    41  jjmod area=2.565     
RS4    47    41               4.406ohm  *SHUNT=11.300
b5    41    43  jjmod area=2.825     
RS5    41    43               3.999ohm  *SHUNT=11.300
b6    48    52  jjmod area=2.170     
RS6    48    52               5.207ohm  *SHUNT=11.300
*FIX
b7    49    42  jjmod area=2.251     
RS7    49    42               5.021ohm  *SHUNT=11.300
b8    42    44  jjmod area=1.471     
RS8    42    44               7.682ohm  *SHUNT=11.300
b9    40    39  jjmod area=1.000     
RS9    40    39              11.300ohm  *SHUNT=11.300
*FIX
b10    32    35  jjmod area=1.523     
RS10    32    35               7.420ohm  *SHUNT=11.300
b11    30    31  jjmod area=2.030     
RS11    30    31               5.567ohm  *SHUNT=11.300
*FIX

XI3              ijtl         16         17
XI5              ijtl         18         19
XI1              ijtl         20         21
XI7               jtl         22          9          4
XI4               jtl         17         23          4
XI6               jtl         19         24          4
XI2               jtl         21         14          4
XI8              sink          9          4

Vindin            20         0  PWL(0ps 0mv 150ps 0mv 151ps 2.068mv 152ps 0mv 250ps 0mv 251ps 2.068mv 252ps 0mv)
Vinclk            18         0  PULSE(0mv 1.034mv 100ps 1ps 1ps 1ps 100ps)
Vinrst            16         0  PWL(0ps 0mv 450ps 0mv 451ps 2.068mv 452ps 0mv 550ps 0mv 551ps 2.068mv 552ps 0mv)
vb     4     0   PWL(0ps 0mV    50ps                  2.500mV)
*FIX
*** netlist file ***

*** jsim input file ***

*** jsim input file ***


.tran 0.1ps 750ps 0ps 0.2ps:
.FILE CIRCUIT108552.CSV


.print phase B2
.print phase B5
.print phase B8
.print phase B11

.end
